`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/18/2020 02:55:21 PM
// Design Name: 
// Module Name: vga_sync
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module vga_sync(
    input  clk    , reset  ,
    input  [11:0] sw,
    output         hsync  , vsync  ,
    output  [ 9:0] pixel_x, pixel_y,
    output  [11:0] rgb
    );
    
    
    
    
    
endmodule    